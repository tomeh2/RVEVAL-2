--===============================================================================
--MIT License

--Copyright (c) 2022 Tomislav Harmina

--Permission is hereby granted, free of charge, to any person obtaining a copy
--of this software and associated documentation files (the "Software"), to deal
--in the Software without restriction, including without limitation the rights
--to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
--copies of the Software, and to permit persons to whom the Software is
--furnished to do so, subject to the following conditions:

--The above copyright notice and this permission notice shall be included in all
--copies or substantial portions of the Software.

--THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
--IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
--FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
--AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
--LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
--OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
--SOFTWARE.
--===============================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use WORK.PKG_CPU.ALL;
use WORK.PKG_FU.ALL;

-- MODULES --
-- 1) ADDRESS GENERATION UNIT
-- 2) STORE DATA

-- Currently both data and address are generated by a single uop. Logic might become more complicated in the future when address calculations for
-- STORE instruction could be fired earlier then data generation

entity execution_unit_1 is
    port(
        cdb : in cdb_type;
        eu_in_0 : in eu_input_type;
    
        valid : in std_logic;       -- Signals that the input values are valid
        ready : out std_logic;      -- Whether this EU is ready to start executing a new operation
        
        -- TO LOAD-STORE UNIT
        lsu_generated_address : out std_logic_vector(CPU_ADDR_WIDTH_BITS - 1 downto 0);
        lsu_generated_data : out std_logic_vector(CPU_DATA_WIDTH_BITS - 1 downto 0);
        lsu_generated_data_tag : out std_logic_vector(PHYS_REGFILE_ADDR_BITS - 1 downto 0);
        lsu_generated_data_valid : out std_logic;
        lsu_stq_tag : out std_logic_vector(STORE_QUEUE_TAG_BITS - 1 downto 0);
        lsu_stq_tag_valid : out std_logic;
        lsu_ldq_tag : out std_logic_vector(LOAD_QUEUE_TAG_BITS - 1 downto 0);
        lsu_ldq_tag_valid : out std_logic;
        
        clk : in std_logic;
        reset : in std_logic
    );
end execution_unit_1;

architecture rtl of execution_unit_1 is
    signal pipeline_reg_0 : exec_unit_1_pipeline_reg_0_type;
    signal pipeline_reg_0_next : exec_unit_1_pipeline_reg_0_type;
    
    alias uop_is_store : std_logic is eu_in_0.operation_select(7);
begin
    process(clk)
    begin
        if (rising_edge(clk)) then
            if (reset = '1') then
                pipeline_reg_0 <= EU_1_PIPELINE_REG_0_INIT;
            else
                pipeline_reg_0 <= pipeline_reg_0_next;
            end if;
        end if;
    end process;
    
    pipeline_reg_0_next.generated_address <= std_logic_vector(unsigned(eu_in_0.operand_2) + unsigned(eu_in_0.immediate)) when eu_in_0.operation_select(6) = '0' else eu_in_0.operand_2;
    pipeline_reg_0_next.generated_data <= eu_in_0.operand_1;
    pipeline_reg_0_next.generated_data_tag <= eu_in_0.phys_src_reg_2_addr;
    pipeline_reg_0_next.generated_data_valid <= uop_is_store and valid;
    pipeline_reg_0_next.ldq_tag <= eu_in_0.ldq_tag;
    pipeline_reg_0_next.ldq_tag_valid <= not uop_is_store and valid;
    pipeline_reg_0_next.stq_tag <= eu_in_0.stq_tag;
    pipeline_reg_0_next.stq_tag_valid <= uop_is_store and valid;
    pipeline_reg_0_next.speculated_branches_mask <= eu_in_0.speculated_branches_mask when cdb.cdb_branch.valid = '0' else eu_in_0.speculated_branches_mask and not cdb.cdb_branch.branch_mask;
    pipeline_reg_0_next.valid <= '1' when valid = '1' and not ((eu_in_0.speculated_branches_mask and cdb.cdb_branch.branch_mask) /= BRANCH_MASK_ZERO and cdb.cdb_branch.branch_mispredicted = '1' and cdb.cdb_branch.valid = '1') else '0';

    lsu_generated_address <= pipeline_reg_0.generated_address;
    lsu_generated_data <= pipeline_reg_0.generated_data;
    lsu_generated_data_tag <= pipeline_reg_0.generated_data_tag;
    lsu_generated_data_valid <= pipeline_reg_0.generated_data_valid and pipeline_reg_0.valid;
    lsu_stq_tag <= pipeline_reg_0.stq_tag;
    lsu_stq_tag_valid <= pipeline_reg_0.stq_tag_valid and pipeline_reg_0.valid;
    lsu_ldq_tag <= pipeline_reg_0.ldq_tag;
    lsu_ldq_tag_valid <= pipeline_reg_0.ldq_tag_valid and pipeline_reg_0.valid;

    ready <= '1';       -- Always ready

end rtl;
